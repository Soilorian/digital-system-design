library verilog;
use verilog.vl_types.all;
entity a is
    port(
        x               : out    vl_logic;
        y               : out    vl_logic
    );
end a;
