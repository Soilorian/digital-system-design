library verilog;
use verilog.vl_types.all;
entity buffer_TB is
end buffer_TB;
