library verilog;
use verilog.vl_types.all;
entity TB_multiplier is
end TB_multiplier;
