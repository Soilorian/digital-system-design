library verilog;
use verilog.vl_types.all;
entity TB_encoder is
end TB_encoder;
